*** LUT Generation for Analog Design ***
.include param130.inc

.include 130nm_NMOS.pm

*** Voltage Sources ***
vdrain	drain 	0	dc 0
Vsource	source  0	dc 0
Vgate	gate	0	dc 0
Vbulk   bulk	0	dc 0

*** Circuit ***
m1	drain gate source bulk nmos w=width l=length ps=p_source pd=p_drain as=a_source ad=a_drain

*** Analysis ***
.save @m1[l]
.save @m1[vgs]
.save @m1[vds]
.save @m1[igd]
.save @m1[igs]
.save @m1[id]
.save @m1[gm]
.save @m1[gmbs]
.save @m1[gds]
.save @m1[cgg]
.save @m1[cgs]
.save @m1[cgd]
.save @m1[cdg]
.save @m1[cgb]
.save @m1[cdd]
.save @m1[csg]

.control
dc vdrain 0 1.3 0.01 vgate 0 1.3 0.01

print @m1[vgs] @m1[vds] @m1[igd] @m1[igs] @m1[id] @m1[gm] @m1[gmbs] @m1[gds] @m1[cgg] @m1[cgs] @m1[cgd] @m1[cdg] @m1[cgb] @m1[cdd] @m1[csg]

.endc

.end
